* eeschema netlist version 1.1 (spice format) creation date: sunday 09 december 2012 04:06:26 pm ist

* Plotting option vplot8_1
r2  2 0 1000
v2  2 0 pwl(0 0 2.6 0 2.60000000001 5 3 5 )
r3  6 0 1000
v3  6 0 pulse(0 5 0 0 0 0.5 1)
r4  1 0 1000
v4  1 0 5
v1  11 0 5
r1  11 0 1000
* 74hc74
a1 [2 6 11 1] [2_in 6_in 11_in 1_in] u1adc
a2 2_in 6_in ~11_in ~1_in 10_out 3_out u1
a3 [10_out 3_out] [10 3]  u1dac
a4 [10 6 11 1] [10_in 6_in 11_in 1_in] u1adc
a5 10_in 6_in ~11_in ~1_in 4_out 5_out u1
a6 [4_out 5_out] [4 5]  u1dac
.model u1 d_dff
.model u1adc adc_bridge(in_low=0.8 in_high=2.0)
.model u1dac dac_bridge(out_low=0.25 out_high=5.0 out_undef=1.8 t_rise=0.5e-9 t_fall=0.5e-9)

.tran  10e-03 4e-00 0e-00
.plot v(6) v(2) v(10) 
.end
