* EESchema Netlist Version 1.1 (Spice format) creation date: Wednesday 15 May 2013 10:41:20 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
v1  6 0 AC		
R3  7 0 R		
U3  7 VPLOT8_1		
C1  7 3 1.59n		
U4  1 3 IPLOT		
U1  5 1 IPLOT		
U2  1 4 IPLOT		
R2  7 4 10000		
R1  5 6 1000		
X1  1 0 7 UA741		

.end
