* EESchema Netlist Version 1.1 (Spice format) creation date: Tuesday 16 April 2013 12:27:13 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
v1  7 0 PULSE		
R1  1 0 5000		
U2  2 7 6 VPLOT8_1		
U1  2 0 IPLOT		
R2  4 5 10000		
U3  5 7 IPLOT		
v2  4 0 10V		
U4  6 1 IPLOT		
Q1  6 2 7 NPN		

.end
