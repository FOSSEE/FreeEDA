* eeschema netlist version 1.1 (spice format) creation date: wednesday 15 may 2013 09:29:30 pm ist
.include ua741.sub

r3  1 7 100k
* Plotting option vplot8_1
V_u1 5 2 0
V_u2 2 3 0
r2  1 3 1000
v1  6 0 10
r1  5 6 10
x1  2 0 7 ua741

.dc  v1 0e-00 5e-00 5e-03
.plot v(1) 
.plot i(V_u1)
.plot i(V_u2)
.end
