* eeschema netlist version 1.1 (spice format) creation date: friday 24 may 2013 02:23:51 pm ist

v1  1 0 sine(0 5 300 0 0)
* Plotting option vplot8_1
r1  3 1 1k
c1  0 3 1u

.tran  5e-03 30e-03 0e-00
.plot v(1) v(3) 
.end
