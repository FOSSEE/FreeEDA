* eeschema netlist version 1.1 (spice format) creation date: monday 13 may 2013 01:31:53 pm ist

V_u3 5 1 0
V_u1 3 8 0
V_u2 1 7 0
v3  4 0 5v
r2  4 2 10000
r1  5 0 1000
v2  0 6 5v
v1  3 0 5v
q2 6 2 7 pnp
q1 8 2 1 npn

.dc  v3 0e-00 5e-00 1e-00
.plot i(V_u3)
.plot i(V_u1)
.plot i(V_u2)
.end
