* eeschema netlist version 1.1 (spice format) creation date: sunday 09 december 2012 03:22:39 pm ist
.include 1n4007.lib

* Plotting option vplot1
* Plotting option vplot
v1  4 1 sine(0 5 50 0 0)
c1  3 0 1e-06
d4  0 1 1n4007
d2  1 3 1n4007
d3  0 4 1n4007
d1  4 3 1n4007
r1  3 0 100000

.tran  100e-06 40e-03 0e-00
.plot v(3)
.plot v(4)-v(1)
.end
