* EESchema Netlist Version 1.1 (Spice format) creation date: Wednesday 15 May 2013 06:59:18 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
U2  4 3 IPLOT		
v1  1 0 DC		
v2  0 5 DC		
U1  3 VPLOT8_1		
Q1  2 0 3 NPN		
R1  1 4 5k		
R2  2 5 7.07k		

.end
