* EESchema Netlist Version 1.1 (Spice format) creation date: Monday 15 April 2013 12:08:03 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
v2  1 0 DC		
U1  3 1 IPLOT		
D1  5 3 DIODE		
R1  2 5 100		
v1  2 0 SINE		

.end
