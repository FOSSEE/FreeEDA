* eeschema netlist version 1.1 (spice format) 
* creation date: thursday 27 september 2012 02:26:44 pm ist

i2  4 0 dc 1
r5  4 0 1
r2  3 1 1
r4  4 3 2
r3  3 0 1
r1  1 0 1
i1  1 0 dc 1
.op
.end

