* EESchema Netlist Version 1.1 (Spice format) creation date: Monday 15 April 2013 10:01:31 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
U2  1 3 7 VPLOT8_1		
R2  1 0 50000		
R1  5 1 100000		
R4  4 0 3000		
U4  7 4 IPLOT		
v1  5 0 15V		
U3  6 3 IPLOT		
R3  5 6 5000		
Q1  7 1 3 NPN		

.end
