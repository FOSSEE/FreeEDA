V1 1 0 dc 1.8
M1 3 1 2 P (20e-6 0.18e-6 -0.4 8.56e-3)
M2 3 0 2 N (10e-6 0.18e-6 0.4 8.56e-3)
V2 2 0 sweep 0 
.dc 0 1.8 0.05
.plot v(3)
.end
