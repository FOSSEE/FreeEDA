* Bridge Rectifier
V1 1 2 sine (5 50)
D1 1 3 mymodel (1e-8 0.026) 
D2 2 3 mymodel (1e-8 0.026)
D3 0 1 mymodel (1e-8 0.026)
D4 0 2 mymodel (1e-8 0.026)
R1 3 0 1
.tran 0.0005 0.04 0
.plot v(1)-v(2) v(3)
.end
