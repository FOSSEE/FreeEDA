* Example to explain modified nodal analyis
V1 1 0 dc 5
R1 1 2 1
R2 2 0 1
R3 2 3 1
R4 1 3 1
V2 3 0 dc 10
.op
.end
