V1 1 0 dc 5
X2 1 2 myR (2)
R3 2 0 1
.op 
.end
