* eeschema netlist version 1.1 (spice format) creation date: thursday 18 april 2013 10:25:46 am ist
.include ua741.sub

v1  5 0 pulse(1 0 0 0 0 0.001 0.002)
c1  6 1 10n
V_u4 2 1 0
* Plotting option vplot8_1
V_u1 4 2 0
V_u2 2 3 0
r2  6 3 1000000
r1  4 5 10000
x1  2 0 6 ua741

.tran  1e-03 2e-03 0e-00
.plot v(5) 
.plot i(V_u4)
.plot v(6) 
.plot i(V_u1)
.plot i(V_u2)
.end
