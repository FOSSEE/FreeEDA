* eeschema netlist version 1.1 (spice format) creation date: monday 13 may 2013 12:54:07 pm ist

* Plotting option vplot8_1
v2  1 0 10v
v1  0 4 10v
V_u1 5 0 0
V_u2 1 7 0
d2  6 3 diode
r2  7 6 5k
r1  4 3 10k
d1  5 3 diode

.dc  v2 0e-00 10e-00 1e-00
.plot v(6) 
.plot i(V_u1)
.plot i(V_u2)
.end
