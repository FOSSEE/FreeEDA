* EESchema Netlist Version 1.1 (Spice format) creation date: Sunday 09 December 2012 04:06:26 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
U2  6 2 10 VPLOT8_1		
R2  2 0 1000		
v2  2 0 PWL		
R3  6 0 1000		
v3  6 0 PULSE		
R4  1 0 1000		
v4  1 0 5		
v1  11 0 5		
R1  11 0 1000		
U1  1 2 6 11 10 3 0 5 4 11 6 10 1 7 74HC74		

.end
