* eeschema netlist version 1.1 (spice format) creation date: monday 13 may 2013 12:59:00 pm ist
.include diode.lib

* Plotting option vplot8_1
V_u2 3 0 0
d1  2 3 diode
r1  1 2 1000
v1  1 0 5v

.dc v1 0e-00 5e-00 50e-03
.plot v(2) 
.plot i(V_u2)
.end
