* EESchema Netlist Version 1.1 (Spice format) creation date: Tuesday 16 April 2013 12:03:45 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
Q1  7 1 5 PNP		
v1  7 0 PULSE		
R1  6 0 5000		
U2  1 7 5 VPLOT8_1		
U1  1 0 IPLOT		
R2  3 4 10000		
U3  4 7 IPLOT		
v2  3 0 10V		
U4  5 6 IPLOT		

.end
