* EESchema Netlist Version 1.1 (Spice format) creation date: Sunday 09 December 2012 08:37:15 AM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
U1  8 4 9 VPLOT8_1		
U12  5 6 9 0 3 74HC86		
U8  8 4 10 0 3 74LS32		
U7  8 4 2 0 3 74LS08		
U9  7 2 10 0 3 74HC02		
U11  7 6 0 3 74HC04		
U10  2 10 5 0 3 7400		
R3  8 0 1000		
v2  8 0 PULSE		
R2  9 0 1000		
R1  4 0 1000		
v1  4 0 PULSE		

.end
