* EESchema Netlist Version 1.1 (Spice format) creation date: Monday 15 April 2013 03:25:12 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
v1  3 0 DC		
U1  0 1 VPLOT8		
R2  1 0 2000		
R1  3 1 500		
D1  0 1 ZENER		

.end
