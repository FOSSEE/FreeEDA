V1 1 0 ac 5
R1 1 2 100
C1 2 0 1e-6 
.ac lin 10 1 10000 
.plot v(2)
.end
