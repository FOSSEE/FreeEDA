V1 1 0 dc 5
R1 1 2 1000
R2 2 3 1000
C1 3 0 0.1e-6 ic=3 
.tran 0 0.5e-3 0.01e-3 UIC 
.ic v(2)=1
.print v(3)
.end
