* eeschema netlist version 1.1 (spice format) creation date: friday 26 april 2013 03:55:55 pm ist
.include npn.lib

i1  5 0 idc
V_u4 0 1 0
V_u2 3 5 0
V_u3 4 6 0
* Plotting option vplot8_1
v1  4 0 2
q1 6 3 1 npn

.dc  v1 0e-00 2e-00 2e-03
.plot i(V_u4)
.plot i(V_u2)
.plot i(V_u3)
.plot v(6) v(1) 
.end
