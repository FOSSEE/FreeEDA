* eeschema netlist version 1.1 (spice format) creation date: wednesday 17 april 2013 12:50:50 pm ist
.include ua741.sub

r3  6 0 1000
v1  5 0 sine(0 5 50 0 0)
* Plotting option vplot8_1
V_u1 4 2 0
V_u2 2 3 0
r2  6 3 9000
r1  4 5 1000
x1  2 0 6 ua741

.tran  10e-03 20e-03 0e-00
.plot v(6) 
.plot i(V_u1)
.plot i(V_u2)
.end
