V1 2 0 dc 0
M1 1 0 2 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
V2 3 0 sweep 0
V3 3 1 dc 0
.dc 0 1.8 0.1
.plot i(V3)
.end
