V1 2 0 dc 2.5
M1 1 0 2 N (20e-6 0.18e-6 1 1e-3 1e-1)
V2 3 0 sweep 0
V3 3 1 dc 0
.dc 0 5 0.1
.plot i(V3)
.end
