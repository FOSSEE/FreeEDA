* eeschema netlist version 1.1 (spice format) creation date: monday 17 december 2012 11:49:47 am ist

* Printing option vprint1
i2  1 0 1
r5  1 0 1
r2  4 3 1
r4  1 4 2
r3  4 0 1
r1  3 0 1
i1  3 0 1

.op
.print v(4)
.end
