* eeschema netlist version 1.1 (spice format) creation date: friday 24 may 2013 01:58:56 pm ist

* Plotting option vplot8_1
v1  1 0 ac 2
r1  3 1 1k
c1  0 3 1u

.ac lin 10 1Hz 10Meg
.plot v(1) v(3) 
.end
