V1 1 0 dc 1.8
M1 3 1 2 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M2 3 0 2 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M3 4 1 3 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M4 4 0 3 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M5 5 1 4 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M6 5 0 4 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M7 6 1 5 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M8 6 0 5 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M9 7 1 6 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M10 7 0 6 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M11 8 1 7 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M12 8 0 7 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M13 9 1 8 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M14 9 0 8 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M15 10 1 9 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M16 10 0 9 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M17 11 1 10 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M18 11 0 10 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M19 12 1 11 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M20 12 0 11 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M21 13 1 12 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M22 13 0 12 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M23 14 1 13 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M24 14 0 13 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M25 15 1 14 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M26 15 0 14 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M27 16 1 15 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M28 16 0 15 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M29 17 1 16 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M30 17 0 16 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M31 18 1 17 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M32 18 0 17 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M33 19 1 18 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M34 19 0 18 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M35 20 1 19 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M36 20 0 19 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M37 21 1 20 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M38 21 0 20 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M39 22 1 21 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M40 22 0 21 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M41 23 1 22 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M42 23 0 22 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M43 24 1 23 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M44 24 0 23 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M45 25 1 24 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M46 25 0 24 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M47 26 1 25 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M48 26 0 25 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M49 27 1 26 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M50 27 0 26 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M51 28 1 27 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M52 28 0 27 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M53 29 1 28 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M54 29 0 28 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M55 30 1 29 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M56 30 0 29 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M57 31 1 30 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M58 31 0 30 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M59 32 1 31 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M60 32 0 31 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
M61 2 1 32 P (20e-6 0.18e-6 -0.4 1e-3 1e-1)
M62 2 0 32 N (20e-6 0.18e-6 0.4 1e-3 1e-1)
.tran 0 20e-9 1e-9
.plot v(2)
.end
