* EESchema Netlist Version 1.1 (Spice format) creation date: Wednesday 15 May 2013 09:29:30 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
R3  1 7 100k		
U3  1 VPLOT8_1		
U1  5 2 IPLOT		
U2  2 3 IPLOT		
R2  1 3 1000		
v1  6 0 10		
R1  5 6 10		
X1  2 0 7 UA741		

.end
