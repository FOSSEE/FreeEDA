* linear circuit
V1 1 0 dc 1
R1 1 2 1
R2 2 0 1
E1 2 3 4 5 0.5
I1 0 3 dc 1
R3 4 0 1
R4 3 4 1
G1 3 5 0 4 0.5
R5 5 4 0.5
R6 5 0 1
.op
.end
