* eeschema netlist version 1.1 (spice format) creation date: tuesday 16 april 2013 11:31:17 am ist

r1  5 7 80000
* Plotting option vplot8_1
r2  7 0 40000
r4  4 0 3300
V_u4 1 4 0
v1  5 0 12v
V_u3 6 2 0
r3  5 6 4000
q1 2 7 1 npn

.dc  v1 0e-00 12e-00 12e-03
.plot v(7) v(2) v(1) 
.plot i(V_u4)
.plot i(V_u3)
.end
