V1 1 0 dc 5
R1 1 2 1e3
C1 2 0 0.1e-6
.tran 0 5e-3 0.5e-3
.plot v(2)
.end
