* EESchema Netlist Version 1.1 (Spice format) creation date: Friday 24 May 2013 01:58:56 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
U1  1 3 VPLOT8_1		
v1  1 0 AC		
R1  3 1 1k		
C1  0 3 1u		

.end
