* EESchema Netlist Version 1.1 (Spice format) creation date: Monday 15 April 2013 08:10:56 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
U3  4 6 VPLOT8_1		
v1  3 5 10		
R2  6 3 2000		
U2  6 2 IPLOT		
U1  4 1 IPLOT		
R1  5 1 1000		
Q1  2 0 4 PNP		

.end
