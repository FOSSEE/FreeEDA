* EESchema Netlist Version 1.1 (Spice format) creation date: Monday 15 April 2013 04:09:24 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
U3  6 7 VPLOT8_1		
U2  7 3 IPLOT		
U1  5 6 IPLOT		
v1  2 0 4		
v2  4 0 10V		
R2  3 0 3300		
R1  4 5 4700		
Q1  7 2 6 NPN		

.end
