* eeschema netlist version 1.1 (spice format) creation date: wednesday 15 may 2013 10:41:20 pm ist
.include ua741.sub

v1  6 0 ac 1
r3  7 0 r
* Plotting option vplot8_1
c1  7 3 1.59n
V_u4 1 3 0
V_u1 5 1 0
V_u2 1 4 0
r2  7 4 10000
r1  5 6 1000
x1  1 0 7 ua741

.ac lin 10 1Hz 1Meg
.plot v(7) 
.plot i(V_u4)
.plot i(V_u1)
.plot i(V_u2)
.end
