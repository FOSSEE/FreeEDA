* EESchema Netlist Version 1.1 (Spice format) creation date: Tuesday 14 May 2013 02:41:09 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
v1  1 0 DC		
U1  5 VPLOT8_1		
U2  4 0 IPLOT		
R2  3 2 20m		
v2  2 4 65m		
R1  1 5 1000		
D1  5 3 DIODE		

.end
