* EESchema Netlist Version 1.1 (Spice format) creation date: Friday 26 April 2013 03:55:55 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
i1  5 0 IDC		
U4  0 1 IPLOT		
U2  3 5 IPLOT		
U3  4 6 IPLOT		
U1  6 1 VPLOT8_1		
v1  4 0 2		
Q1  1 3 6 NPN		

.end
