* eeschema netlist version 1.1 (spice format) creation date: monday 17 december 2012 11:47:07 am ist

* Printing option vprint1
r3  2 4 1
r4  2 3 1
r1  4 3 1
r2  4 0 1
v2  2 0 10
v1  3 0 5

.op
.print v(4)
.end
